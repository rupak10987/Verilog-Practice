`timescale 1ns/1ps
module comb1_tb();